`ifndef CONSTANT
// ALU operations {inst [30], funct3}
`define ALU_ADD                 3'b001
`define ALU_SUB                 3'b010
`define ALU_MULT                3'b011
`define ALU_INV                 3'b100
`define ALU_NOP                 3'b000

`endif
